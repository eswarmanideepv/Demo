// example.v
module main;
    initial begin
        $display("Hello, Icarus Verilog!");
        $display("Manideep");
        $finish;
    end
endmodule